`define MPF_DISABLED 1
